netcdf drydep_tables {
dimensions:
  n_species_table = 192;
  NHen  = 6;
  chars = 16;
variables:
  
  char species_name_table(n_species_table,chars);
    species_name_table:long_name = "names of species in dry deposition tables" ;
  double dfoxd(n_species_table);
    dfoxd:long_name = "data for foxd (reactivity factor for oxidation)";
  double dheff(n_species_table,NHen);
    dheff:long_name = "data for effective Henry's Law coefficient";
  double mol_wghts(n_species_table);
    mol_wghts:long_name = "species molecular mass";
    mol_wghts:units = "grams/mole";
    
// global attributes:

  :Created_by = "Francis Vitt";
  :Source = "Data extracted from cime source code src/drivers/mct/shr/seq_drydep_mod.F90, tag cime5.8.26";

data:

  species_name_table =
         "OX              ",
         "H2O2            ",
         "OH              ",
         "HO2             ",
         "CO              ",
         "CH4             ",
         "CH3O2           ",
         "CH3OOH          ",
         "CH2O            ",
         "HCOOH           ",
         "NO              ",
         "NO2             ",
         "HNO3            ",
         "CO2             ",
         "NH3             ",
         "N2O5            ",
         "NO3             ",
         "CH3OH           ",
         "HO2NO2          ",
         "O1D             ",
         "C2H6            ",
         "C2H5O2          ",
         "PO2             ",
         "MACRO2          ",
         "ISOPO2          ",
         "C4H10           ",
         "CH3CHO          ",
         "C2H5OOH         ",
         "C3H6            ",
         "POOH            ",
         "C2H4            ",
         "PAN             ",
         "CH3COOOH        ",
         "MTERP           ",
         "GLYOXAL         ",
         "CH3COCHO        ",
         "GLYALD          ",
         "CH3CO3          ",
         "C3H8            ",
         "C3H7O2          ",
         "CH3COCH3        ",
         "C3H7OOH         ",
         "RO2             ",
         "ROOH            ",
         "Rn              ",
         "ISOP            ",
         "MVK             ",
         "MACR            ",
         "C2H5OH          ",
         "ONITR           ",
         "ONIT            ",
         "ISOPNO3         ",
         "HYDRALD         ",
         "HCN             ",
         "CH3CN           ",
         "SO2             ",
         "SOAGff0         ",
         "SOAGff1         ",
         "SOAGff2         ",
         "SOAGff3         ",
         "SOAGff4         ",
         "SOAGbg0         ",
         "SOAGbg1         ",
         "SOAGbg2         ",
         "SOAGbg3         ",
         "SOAGbg4         ",
         "SOAG0           ",
         "SOAG1           ",
         "SOAG2           ",
         "SOAG3           ",
         "SOAG4           ",
         "IVOC            ",
         "SVOC            ",
         "IVOCbb          ",
         "IVOCff          ",
         "SVOCbb          ",
         "SVOCff          ",
         "N2O             ",
         "H2              ",
         "C2H2            ",
         "CH3COOH         ",
         "EOOH            ",
         "HYAC            ",
         "BIGENE          ",
         "BIGALK          ",
         "MEK             ",
         "MEKOOH          ",
         "MACROOH         ",
         "MPAN            ",
         "ALKNIT          ",
         "NOA             ",
         "ISOPNITA        ",
         "ISOPNITB        ",
         "ISOPNOOH        ",
         "NC4CHO          ",
         "NC4CH2OH        ",
         "TERPNIT         ",
         "NTERPOOH        ",
         "ALKOOH          ",
         "BIGALD          ",
         "HPALD           ",
         "IEPOX           ",
         "XOOH            ",
         "ISOPOOH         ",
         "TOLUENE         ",
         "CRESOL          ",
         "TOLOOH          ",
         "BENZENE         ",
         "PHENOL          ",
         "BEPOMUC         ",
         "PHENOOH         ",
         "C6H5OOH         ",
         "BENZOOH         ",
         "BIGALD1         ",
         "BIGALD2         ",
         "BIGALD3         ",
         "BIGALD4         ",
         "TEPOMUC         ",
         "BZOOH           ",
         "BZALD           ",
         "PBZNIT          ",
         "XYLENES         ",
         "XYLOL           ",
         "XYLOLOOH        ",
         "XYLENOOH        ",
         "BCARY           ",
         "TERPOOH         ",
         "TERPROD1        ",
         "TERPROD2        ",
         "TERP2OOH        ",
         "DMS             ",
         "H2SO4           ",
         "HONITR          ",
         "MACRN           ",
         "MVKN            ",
         "ISOPN2B         ",
         "ISOPN3B         ",
         "ISOPN4D         ",
         "ISOPN1D         ",
         "ISOPNOOHD       ",
         "ISOPNOOHB       ",
         "ISOPNBNO3       ",
         "NO3CH2CHO       ",
         "HYPERACET       ",
         "HCOCH2OOH       ",
         "DHPMPAL         ",
         "MVKOOH          ",
         "ISOPOH          ",
         "ISOPFDN         ",
         "ISOPFNP         ",
         "INHEB           ",
         "HMHP            ",
         "HPALD1          ",
         "INHED           ",
         "HPALD4          ",
         "ISOPHFP         ",
         "HPALDB1C        ",
         "HPALDB4C        ",
         "ICHE            ",
         "ISOPFDNC        ",
         "ISOPFNC         ",
         "TERPNT          ",
         "TERPNS          ",
         "TERPNT1         ",
         "TERPNS1         ",
         "TERPNPT         ",
         "TERPNPS         ",
         "TERPNPT1        ",
         "TERPNPS1        ",
         "TERPFDN         ",
         "SQTN            ",
         "TERPHFN         ",
         "TERP1OOH        ",
         "TERPDHDP        ",
         "TERPF2          ",
         "TERPF1          ",
         "TERPA           ",
         "TERPA2          ",
         "TERPK           ",
         "TERPAPAN        ",
         "TERPACID        ",
         "TERPA2PAN       ",
         "APIN            ",
         "BPIN            ",
         "LIMON           ",
         "MYRC            ",
         "TERPACID2       ",
         "TERPACID3       ",
         "TERPA3PAN       ",
         "TERPOOHL        ",
         "TERPA3          ",
         "TERP2AOOH       " ;

  dfoxd = 
        1.       // OX
       ,1.       // H2O2
       ,1.       // OH
       ,.1       // HO2
       ,1.e-36   // CO
       ,1.e-36   // CH4
       ,1.       // CH3O2
       ,1.       // CH3OOH
       ,1.       // CH2O
       ,1.       // HCOOH
       ,0.       // NO
       ,.1       // NO2
       ,1.e-36   // HNO3
       ,1.e-36   // CO2
       ,1.e-36   // NH3
       ,.1       // N2O5
       ,1.       // NO3
       ,1.       // CH3OH
       ,.1       // HO2NO2
       ,1.       // O1D
       ,1.e-36   // C2H6
       ,.1       // C2H5O2
       ,.1       // PO2
       ,.1       // MACRO2
       ,.1       // ISOPO2
       ,1.e-36   // C4H10
       ,1.       // CH3CHO
       ,1.       // C2H5OOH
       ,1.e-36   // C3H6
       ,1.       // POOH
       ,1.e-36   // C2H4
       ,.1       // PAN
       ,1.       // CH3COOOH
       ,1.e-36   // MTERP
       ,1.       // GLYOXAL
       ,1.       // CH3COCHO
       ,1.       // GLYALD
       ,.1       // CH3CO3
       ,1.e-36   // C3H8
       ,.1       // C3H7O2
       ,1.       // CH3COCH3
       ,1.       // C3H7OOH
       ,.1       // RO2
       ,1.       // ROOH
       ,1.e-36   // Rn
       ,1.e-36   // ISOP
       ,1.       // MVK
       ,1.       // MACR
       ,1.       // C2H5OH 
       ,1.       // ONITR
       ,.1       // ONIT
       ,.1       // ISOPNO3
       ,1.       // HYDRALD
       ,1.e-36   // HCN
       ,1.e-36   // CH3CN
       ,1.e-36   // SO2
       ,0.1      // SOAGff0
       ,0.1      // SOAGff1
       ,0.1      // SOAGff2
       ,0.1      // SOAGff3
       ,0.1      // SOAGff4
       ,0.1      // SOAGbg0
       ,0.1      // SOAGbg1
       ,0.1      // SOAGbg2
       ,0.1      // SOAGbg3
       ,0.1      // SOAGbg4
       ,0.1      // SOAG0
       ,0.1      // SOAG1
       ,0.1      // SOAG2
       ,0.1      // SOAG3
       ,0.1      // SOAG4
       ,0.1      // IVOC
       ,0.1      // SVOC 
       ,0.1      // IVOCbb
       ,0.1      // IVOCff
       ,0.1      // SVOCbb
       ,0.1      // SVOCff
       ,1.e-36   // N2O
       ,1.e-36   // H2
       ,1.e-36   // C2H2
       ,1.       // CH3COOH
       ,1.       // EOOH
       ,1.       // HYAC
       ,1.e-36   // BIGENE
       ,1.e-36   // BIGALK
       ,1.       // MEK
       ,1.       // MEKOOH
       ,1.       // MACROOH
       ,1.       // MPAN
       ,1.       // ALKNIT
       ,1.       // NOA
       ,1.       // ISOPNITA
       ,1.       // ISOPNITB
       ,1.       // ISOPNOOH
       ,1.       // NC4CHO
       ,1.       // NC4CH2OH
       ,1.       // TERPNIT
       ,1.       // NTERPOOH
       ,1.       // ALKOOH
       ,1.       // BIGALD
       ,1.       // HPALD
       ,1.       // IEPOX
       ,1.       // XOOH
       ,1.       // ISOPOOH
       ,1.e-36   // TOLUENE
       ,1.       // CRESOL
       ,1.       // TOLOOH
       ,1.e-36   // BENZENE
       ,1.       // PHENOL
       ,1.       // BEPOMUC
       ,1.       // PHENOOH
       ,1.       // C6H5OOH
       ,1.       // BENZOOH
       ,1.       // BIGALD1
       ,1.       // BIGALD2
       ,1.       // BIGALD3
       ,1.       // BIGALD4
       ,1.       // TEPOMUC
       ,1.       // BZOOH
       ,1.       // BZALD
       ,1.       // PBZNIT
       ,1.e-36   // XYLENES
       ,1.       // XYLOL
       ,1.       // XYLOLOOH
       ,1.       // XYLENOOH
       ,1.e-36   // BCARY
       ,1.       // TERPOOH
       ,1.       // TERPROD1
       ,1.       // TERPROD2
       ,1.       // TERP2OOH
       ,1.e-36   // DMS
       ,1.e-36   // H2SO4
       ,1.       // HONITR
       ,1.       // MACRN   
       ,1.       // MVKN
       ,1.       // ISOPN2B
       ,1.       // ISOPN3B
       ,1.       // ISOPN4D
       ,1.       // ISOPN1D
       ,1.       // ISOPNOOHD
       ,1.       // ISOPNOOHB
       ,1.       // ISOPNBNO3
       ,1.       // NO3CH2CHO
       ,1.       // HYPERACET
       ,1.       // HCOCH2OOH
       ,1.       // DHPMPAL
       ,1.       // MVKOOH
       ,1.       // ISOPOH
       ,1.       // ISOPFDN
       ,1.       // ISOPFNP
       ,1.       // INHEB
       ,1.       // HMHP
       ,1.       // HPALD1
       ,1.       // INHED
       ,1.       // HPALD4  
       ,1.       // ISOPHFP
       ,1.       // HPALDB1C
       ,1.       // HPALDB4C
       ,1.       // ICHE
       ,1.       // ISOPFDNC
       ,1.       // ISOPFNC
       ,1.       // TERPNT
       ,1.       // TERPNS
       ,1.       // TERPNT1
       ,1.       // TERPNS1
       ,1.       // TERPNPT
       ,1.       // TERPNPS
       ,1.       // TERPNPT1
       ,1.       // TERPNPS1
       ,1.       // TERPFDN
       ,1.       // SQTN
       ,1.       // TERPHFN 
       ,1.       // TERP1OOH
       ,1.       // TERPDHDP
       ,1.       // TERPF2
       ,1.       // TERPF1
       ,1.       // TERPA
       ,1.       // TERPA2 
       ,1.       // TERPK
       ,1.       // TERPAPAN
       ,1.       // TERPACID
       ,1.       // TERPA2PAN
       ,1.e-36   // APIN
       ,1.e-36   // BPIN
       ,1.e-36   // LIMON
       ,1.e-36   // MYRC
       ,1.       // TERPACID2
       ,1.       // TERPACID3
       ,1.       // TERPA3PAN
       ,1.       // TERPOOHL
       ,1.       // TERPA3
       ,1.   ;   // TERP2AOOH

 dheff = 
        1.03e-02, 2830.,  0.,            0., 0.,         0., // OX
        8.70e+04, 7320.,  2.2e-12,   -3730., 0.,         0., // H2O2
        3.90e+01, 4300.,  0.,            0., 0.,         0., // OH
        6.90e+02, 5900.,  0.,            0., 0.,         0., // HO2
        9.81e-04, 1650.,  0.,            0., 0.,         0., // CO
        1.41e-03, 1820.,  0.,            0., 0.,         0., // CH4
        2.38e+00, 5280.,  0.,            0., 0.,         0., // CH3O2
        3.00e+02, 5280.,  0.,            0., 0.,         0., // CH3OOH
        3.23e+03, 7100.,  0.,            0., 0.,         0., // CH2O
        8.90e+03, 6100.,  1.8e-04,     -20., 0.,         0., // HCOOH
        1.92e-03, 1762.,  0.,            0., 0.,         0., // NO
        1.20e-02, 2440.,  0.,            0., 0.,         0., // NO2
        2.10e+05, 8700.,  2.2e+01,       0., 0.,         0., // HNO3
        3.44e-02, 2715.,  4.3e-07,   -1000., 4.7e-11,-1760., // CO2
        6.02e+01, 4160.,  1.7e-05,   -4325., 1.0e-14,-6716., // NH3
        2.14e+00, 3362.,  0.,            0., 0.,         0., // N2O5
        3.80e-02,    0.,  0.,            0., 0.,         0., // NO3
        2.03e+02, 5645.,  0.,            0., 0.,         0., // CH3OH
        4.00e+01, 8400.,  1.3e-06,       0., 0.,         0., // HO2NO2
        1.00e-16,    0.,  0.,            0., 0.,         0., // O1D
        1.88e-03, 2750.,  0.,            0., 0.,         0., // C2H6
        2.38e+00, 5280.,  0.,            0., 0.,         0., // C2H5O2
        2.38e+00, 5280.,  0.,            0., 0.,         0., // PO2
        2.38e+00, 5280.,  0.,            0., 0.,         0., // MACRO2
        2.38e+00, 5280.,  0.,            0., 0.,         0., // ISOPO2
        1.70e-03,    0.,  0.,            0., 0.,         0., // C4H10
        1.29e+01, 5890.,  0.,            0., 0.,         0., // CH3CHO
        3.36e+02, 5995.,  0.,            0., 0.,         0., // C2H5OOH
        5.57e-03, 2800.,  0.,            0., 0.,         0., // C3H6
        1.50e+06, 6014.,  0.,            0., 0.,         0., // POOH
        5.96e-03, 2200.,  0.,            0., 0.,         0., // C2H4
        2.80e+00, 5730.,  0.,            0., 0.,         0., // PAN
        8.37e+02, 5310.,  1.8e-04,     -20., 0.,         0., // CH3COOOH
        2.94e-02, 1800.,  0.,            0., 0.,         0., // MTERP
        4.19e+05, 7480.,  0.,            0., 0.,         0., // GLYOXAL
        3.50e+03, 7545.,  0.,            0., 0.,         0., // CH3COCHO
        4.00e+04, 4630.,  0.,            0., 0.,         0., // GLYALD
        1.00e-01,    0.,  0.,            0., 0.,         0., // CH3CO3
        1.51e-03, 3120.,  0.,            0., 0.,         0., // C3H8
        2.38e+00, 5280.,  0.,            0., 0.,         0., // C3H7O2
        2.78e+01, 5530.,  0.,            0., 0.,         0., // CH3COCH3
        3.36e+02, 5995.,  0.,            0., 0.,         0., // C3H7OOH
        2.38e+00, 5280.,  0.,            0., 0.,         0., // RO2
        3.36e+02, 5995.,  0.,            0., 0.,         0., // ROOH
        0.00e+00,    0.,  0.,            0., 0.,         0., // Rn
        3.45e-02, 4400.,  0.,            0., 0.,         0., // ISOP
        4.10e+01, 6014.,  0.,            0., 0.,         0., // MVK
        6.50e+00, 6014.,  0.,            0., 0.,         0., // MACR
        1.90e+02, 6500.,  0.,            0., 0.,         0., // C2H5OH
        1.44e+03, 6014.,  0.,            0., 0.,         0., // ONITR
        1.00e+03, 6000.,  0.,            0., 0.,         0., // ONIT
        2.38e+00, 5280.,  0.,            0., 0.,         0., // ISOPNO3
        1.10e+05, 6000.,  0.,            0., 0.,         0., // HYDRALD
        9.02e+00, 8258.,  0.,            0., 0.,         0., // HCN
        5.28e+01, 3970.,  0.,            0., 0.,         0., // CH3CN
        1.36e+00, 3100.,  1.30e-02,   1960., 6.6e-08, 1500., // SO2
        1.3e+07,     0.,  0.,            0., 0.,         0., // SOAGff0
        3.2e+05,     0.,  0.,            0., 0.,         0., // SOAGff1
        4.0e+05,     0.,  0.,            0., 0.,         0., // SOAGff2 
        1.3e+05,     0.,  0.,            0., 0.,         0., // SOAGff3
        1.6e+05,     0.,  0.,            0., 0.,         0., // SOAGff4
        7.9e+11,     0.,  0.,            0., 0.,         0., // SOAGbg0
        6.3e+10,     0.,  0.,            0., 0.,         0., // SOAGbg1
        3.2e+09,     0.,  0.,            0., 0.,         0., // SOAGbg2
        6.3e+08,     0.,  0.,            0., 0.,         0., // SOAGbg3
        3.2e+07,     0.,  0.,            0., 0.,         0., // SOAGbg4
        4.0e+11,     0.,  0.,            0., 0.,         0., // SOAG0
        3.2e+10,     0.,  0.,            0., 0.,         0., // SOAG1
        1.6e+09,     0.,  0.,            0., 0.,         0., // SOAG2
        3.2e+08,     0.,  0.,            0., 0.,         0., // SOAG3
        1.6e+07,     0.,  0.,            0., 0.,         0., // SOAG4
        1.e+03,      0.,  0.,            0., 0.,         0., // IVOC
        1.e+03,      0.,  0.,            0., 0.,         0., // SVOC
        1.e+03,      0.,  0.,            0., 0.,         0., // IVOCbb
        1.e+03,      0.,  0.,            0., 0.,         0., // IVOCff
        1.e+03,      0.,  0.,            0., 0.,         0., // SVOCbb
        1.e+03,      0.,  0.,            0., 0.,         0., // SVOCff
        2.42e-02, 2710.,  0.,            0., 0.,         0., // N2O
        7.9e-04,   530.,  0.,            0., 0.,         0., // H2
        4.14e-02, 1890.,  0.,            0., 0.,         0., // C2H2
        4.1e+03,  6200.,  0.,            0., 0.,         0., // CH3COOH
        1.9e+06,  6014.,  0.,            0., 0.,         0., // EOOH
        1.46e+03, 6014.,  0.,            0., 0.,         0., // HYAC
        5.96e-03, 2365.,  0.,            0., 0.,         0., // BIGENE
        1.24e-03, 3010.,  0.,            0., 0.,         0., // BIGALK
        1.80e+01, 5740.,  0.,            0., 0.,         0., // MEK
        6.4e+04,  6014.,  0.,            0., 0.,         0., // MEKOOH
        4.4e+06,  6014.,  0.,            0., 0.,         0., // MACROOH
        1.72e+00, 5700.,  0.,            0., 0.,         0., // MPAN
        1.01e+00, 5790.,  0.,            0., 0.,         0., // ALKNIT
        1.e+03,   6014.,  0.,            0., 0.,         0., // NOA
        8.34e+03, 6014.,  0.,            0., 0.,         0., // ISOPNITA
        4.82e+04, 6014.,  0.,            0., 0.,         0., // ISOPNITB
        8.75e+04, 6014.,  0.,            0., 0.,         0., // ISOPNOOH
        1.46e+03, 6014.,  0.,            0., 0.,         0., // NC4CHO
        4.02e+04, 9500.,  0.,            0., 0.,         0., // NC4CH2OH
        8.41e+03, 6014.,  0.,            0., 0.,         0., // TERPNIT
        6.67e+04, 6014.,  0.,            0., 0.,         0., // NTERPOOH
        3.36e+02, 5995.,  0.,            0., 0.,         0., // ALKOOH
        9.6e+00,  6220.,  0.,            0., 0.,         0., // BIGALD
        2.30e+05, 6014.,  0.,            0., 0.,         0., // HPALD
        3.e+07,   6014.,  0.,            0., 0.,         0., // IEPOX
        1.e+11,   5995.,  0.,            0., 0.,         0., // XOOH
        3.5e+06,  5995.,  0.,            0., 0.,         0., // ISOPOOH
        1.5e-01,  4300.,  0.,            0., 0.,         0., // TOLUENE
        5.67e+02, 5800.,  0.,            0., 0.,         0., // CRESOL
        2.30e+04, 5995.,  0.,            0., 0.,         0., // TOLOOH
        1.8e-01,  3800.,  0.,            0., 0.,         0., // BENZENE
        2.84e+03, 2700.,  0.,            0., 0.,         0., // PHENOL
        3.e+07,   6014.,  0.,            0., 0.,         0., // BEPOMUC
        1.5e+06,  5995.,  0.,            0., 0.,         0., // PHENOOH
        3.36e+02, 5995.,  0.,            0., 0.,         0., // C6H5OOH
        2.3e+03,  5995.,  0.,            0., 0.,         0., // BENZOOH 
        1.e+05,   5890.,  0.,            0., 0.,         0., // BIGALD1 
        2.9e+04,  5890.,  0.,            0., 0.,         0., // BIGALD2
        2.2e+04,  5890.,  0.,            0., 0.,         0., // BIGALD3
        2.2e+04,  5890.,  0.,            0., 0.,         0., // BIGALD4
        2.5e+05,  6014.,  0.,            0., 0.,         0., // TEPOMUC
        3.36e+02, 5995.,  0.,            0., 0.,         0., // BZOOH
        3.24e+01, 6300.,  0.,            0., 0.,         0., // BZALD
        2.8e+00,  5730.,  0.,            0., 0.,         0., // PBZNIT
        2.e-01,   4300.,  0.,            0., 0.,         0., // XYLENES
        1.01e+03, 6800.,  0.,            0., 0.,         0., // XYLOL
        1.9e+06,  5995.,  0.,            0., 0.,         0., // XYLOLOOH
        3.36e+02, 5995.,  0.,            0., 0.,         0., // XYLENOOH
        5.57e-03, 2800.,  0.,            0., 0.,         0., // BCARY
        3.6e+06,  6014.,  0.,            0., 0.,         0., // TERPOOH
        3.92e+04, 6014.,  0.,            0., 0.,         0., // TERPROD1
        7.20e+04, 6014.,  0.,            0., 0.,         0., // TERPROD2
        3.36e+02, 5995.,  0.,            0., 0.,         0., // TERP2OOH
        5.4e-01,  3460.,  0.,            0., 0.,         0., // DMS
        1.e+11,   6014.,  0.,            0., 0.,         0., // H2SO4
        2.64e+03, 6014.,  0.,            0., 0.,         0., // HONITR
        4.14e+06, 6014.,  0.,            0., 0.,         0., // MACRN
        1.84e+05, 6014.,  0.,            0., 0.,         0., // MVKN
        8.34e+03, 6014.,  0.,            0., 0.,         0., // ISOPN2B
        8.34e+03, 6014.,  0.,            0., 0.,         0., // ISOPN3B
        4.82e+04, 6014.,  0.,            0., 0.,         0., // ISOPN4D
        4.82e+04, 6014.,  0.,            0., 0.,         0., // ISOPN1D
        9.67e+04, 6014.,  0.,            0., 0.,         0., // ISOPNOOHD
        6.61e+04, 6014.,  0.,            0., 0.,         0., // ISOPNOOHB
        8.34e+03, 6014.,  0.,            0., 0.,         0., // ISOPNBNO3
        3.39e+04, 6014.,  0.,            0., 0.,         0., // NO3CH2CHO
        1.16e+04, 6014.,  0.,            0., 0.,         0., // HYPERACET
        2.99e+04, 6014.,  0.,            0., 0.,         0., // HCOCH2OOH
        9.37e+07, 6014.,  0.,            0., 0.,         0., // DHPMPAL
        1.24e+06, 6014.,  0.,            0., 0.,         0., // MVKOOH
        8.77e+06, 6014.,  0.,            0., 0.,         0., // ISOPOH
        5.02e+08, 6014.,  0.,            0., 0.,         0., // ISOPFDN
        2.97e+11, 6014.,  0.,            0., 0.,         0., // ISOPFNP
        1.05e+05, 6014.,  0.,            0., 0.,         0., // INHEB
        1.70e+06, 9870.,  0.,            0., 0.,         0., // HMHP
        2.30e+05, 6014.,  0.,            0., 0.,         0., // HPALD1  
        1.51e+05, 6014.,  0.,            0., 0.,         0., // INHED
        2.30e+05, 6014.,  0.,            0., 0.,         0., // HPALD4
        7.60e+09, 6014.,  0.,            0., 0.,         0., // ISOPHFP 
        5.43e+04, 6014.,  0.,            0., 0.,         0., // HPALDB1C
        5.43e+04, 6014.,  0.,            0., 0.,         0., // HPALDB4C
        2.09e+06, 6014.,  0.,            0., 0.,         0., // ICHE
        7.16e+09, 6014.,  0.,            0., 0.,         0., // ISOPFDNC
        1.41e+11, 6014.,  0.,            0., 0.,         0., // ISOPFNC
        8.41e+03, 6014.,  0.,            0., 0.,         0., // TERPNT
        8.41e+03, 6014.,  0.,            0., 0.,         0., // TERPNS
        8.55e+03, 6014.,  0.,            0., 0.,         0., // TERPNT1
        8.55e+03, 6014.,  0.,            0., 0.,         0., // TERPNS1
        6.67e+04, 6014.,  0.,            0., 0.,         0., // TERPNPT
        6.67e+04, 6014.,  0.,            0., 0.,         0., // TERPNPS
        6.78e+04, 6014.,  0.,            0., 0.,         0., // TERPNPT1
        6.78e+04, 6014.,  0.,            0., 0.,         0., // TERPNPS1
        1.65e+09, 6014.,  0.,            0., 0.,         0., // TERPFDN
        9.04e+03, 6014.,  0.,            0., 0.,         0., // SQTN
        7.53e+11, 6014.,  0.,            0., 0.,         0., // TERPHFN
        3.64e+06, 6014.,  0.,            0., 0.,         0., // TERP1OOH
        3.41e+14, 6014.,  0.,            0., 0.,         0., // TERPDHDP
        6.54e+01, 6014.,  0.,            0., 0.,         0., // TERPF2
        4.05e+04, 6014.,  0.,            0., 0.,         0., // TERPF1
        3.92e+04, 6014.,  0.,            0., 0.,         0., // TERPA
        7.20e+04, 6014.,  0.,            0., 0.,         0., // TERPA2
        6.39e+01, 6014.,  0.,            0., 0.,         0., // TERPK
        7.94e+03, 6014.,  0.,            0., 0.,         0., // TERPAPAN
        5.63e+06, 6014.,  0.,            0., 0.,         0., // TERPACID
        9.59e+03, 6014.,  0.,            0., 0.,         0., // TERPA2PAN
        2.94e-02, 1800.,  0.,            0., 0.,         0., // APIN
        1.52e-02, 4500.,  0.,            0., 0.,         0., // BPIN
        4.86e-02, 4600.,  0.,            0., 0.,         0., // LIMON
        7.30e-02, 2800.,  0.,            0., 0.,         0., // MYRC
        2.64e+06, 6014.,  0.,            0., 0.,         0., // TERPACID2
        3.38e+09, 6014.,  0.,            0., 0.,         0., // TERPACID3
        1.23e+07, 6014.,  0.,            0., 0.,         0., // TERPA3PAN
        4.41e+12, 6014.,  0.,            0., 0.,         0., // TERPOOHL
        1.04e+08, 6014.,  0.,            0., 0.,         0., // TERPA3
        3.67e+06, 6014.,  0.,            0., 0.,         0.; // TERP2AOOH

  mol_wghts =
       47.9981995, 34.0135994, 17.0067997, 33.0061989, 28.0104008,
       16.0405998, 47.0320015, 48.0393982, 30.0251999, 46.0246010,
       30.0061398, 46.0055389, 63.0123405, 44.0098000, 17.0289402,
       108.010483, 62.0049400, 32.0400009, 79.0117416, 15.9994001,
       30.0664005, 61.0578003, 91.0830002, 119.093399, 117.119797,
       58.1180000, 44.0509987, 62.0652008, 42.0774002, 92.0904007,
       28.0515995, 121.047943, 76.0497971, 136.228394, 58.0355988,
       72.0614014, 60.0503998, 75.0423965, 44.0922012, 75.0836029,
       58.0768013, 76.0910034, 89.070126,  90.078067,  222.000000,
       68.1141968, 70.0877991, 70.0877991, 46.0657997, 147.125946,
       119.074341, 162.117935, 100.112999, 27.0256,     41.0524,
       64.064800,  250.,       250.,       250.,       250.,      
       250.,       250.,       250.,       250.,       250.,      
       250.,       250.,       250.,       250.,       250.,      
       250.,       170.3,      170.3,      170.3,       170.3,    
       170.3,      170.3,      44.0129,    2.0148,     26.0368,   
       60.0504,    78.0646,    74.0762,    56.1032,    72.1438,   
       72.1026,    104.101,    120.101,    147.085,    133.141,   
       119.074,    147.126,    147.126,    163.125,    145.111,   
       147.126,    215.24,     231.24,     104.143,    98.0982,   
       116.112,    118.127,    150.126,    118.127,    92.1362,   
       108.136,    174.148,    78.1104,    94.1098,    126.109,   
       176.122,    110.109,    160.122,    84.0724,    98.0982,   
       98.0982,    112.124,    140.134,    124.135,    106.121,   
       183.118,    106.162,    122.161,    204.173,    188.174,   
       204.343,    186.241,    168.227,    154.201,    200.226,   
       62.1324,    98.0784,    135.118733, 149.102257, 149.102257,
       147.129469, 147.129469, 147.129469, 147.129469, 163.128874,
       163.128874, 147.129469, 105.049617, 90.078067,  76.05145,  
       136.103494, 120.104089, 102.131897, 226.141733, 197.143565,
       163.128874, 64.040714,  116.11542,  163.128874, 116.11542, 
       150.130112, 116.11542,  116.11542,  116.11542,  224.125851,
       195.127684, 215.246675, 215.246675, 215.246675, 215.246675,
       231.24608,  231.24608,  231.24608,  231.24608,  294.258938,
       283.36388,  265.260771, 186.248507, 236.262604, 110.153964,
       168.233221, 168.233221, 154.206603, 138.207199, 245.229603,
       200.232031, 231.202986, 136.228394, 136.228394, 136.228394,
       136.228394, 186.205413, 202.204818, 247.202391, 218.247317,
       170.206008, 186.248507 ;

}